module or_gate(Y,a,b);
output Y;
input a,b;
or a_1(Y,a,b);
endmodule
