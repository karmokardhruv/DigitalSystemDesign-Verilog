module not_data(a,Y);
input a;
output Y;
assign Y=~a;
endmodule