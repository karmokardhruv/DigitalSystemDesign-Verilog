module xor_gate(Y,a,b);
output Y;
input a, b;
xor a_1(Y,a,b);
endmodule
