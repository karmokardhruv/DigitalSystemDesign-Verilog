module not_gates(Y, a);
output Y; 
input a; 
not a_1(Y,a); 
endmodule