module dec5x32 (
input[4:0]a,
output[31:0]y);
assign y[0] = (~a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0]);
assign y[1] = (~a[4])&(~a[3])&(~a[2])&(~a[1])&(a[0]);
assign y[2] = (~a[4])&(~a[3])&(~a[2])&(a[1])&(~a[0]);
assign y[3] = (~a[4])&(~a[3])&(~a[2])&(a[1])&(a[0]);
assign y[4] = (~a[4])&(~a[3])&(a[2])&(~a[1])&(~a[0]);
assign y[5] = (~a[4])&(~a[3])&(a[2])&(~a[1])&(a[0]);
assign y[6] = (~a[4])&(~a[3])&(a[2])&(a[1])&(~a[0]);
assign y[7] = (~a[4])&(~a[3])&(a[2])&(a[1])&(a[0]);
assign y[8] = (~a[4])&(a[3])&(~a[2])&(~a[1])&(~a[0]);
assign y[9] = (~a[4])&(a[3])&(~a[2])&(~a[1])&(a[0]);
assign y[10] = (~a[4])&(a[3])&(~a[2])&(a[1])&(~a[0]);
assign y[11] = (~a[4])&(a[3])&(~a[2])&(a[1])&(a[0]);
assign y[12] = (~a[4])&(a[3])&(a[2])&(~a[1])&(~a[0]);
assign y[13] = (~a[4])&(a[3])&(a[2])&(~a[1])&(a[0]);
assign y[14] = (~a[4])&(a[3])&(a[2])&(a[1])&(~a[0]);
assign y[15] = (~a[4])&(a[3])&(a[2])&(a[1])&(a[0]);
assign y[16] = (a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0]);
assign y[17] = (a[4])&(~a[3])&(~a[2])&(~a[1])&(a[0]);
assign y[18] = (a[4])&(~a[3])&(~a[2])&(a[1])&(~a[0]);
assign y[19] = (a[4])&(~a[3])&(~a[2])&(a[1])&(a[0]);
assign y[20] = (a[4])&(~a[3])&(a[2])&(~a[1])&(~a[0]);
assign y[21] = (a[4])&(~a[3])&(a[2])&(~a[1])&(a[0]);
assign y[22] = (a[4])&(~a[3])&(a[2])&(a[1])&(~a[0]);
assign y[23] = (a[4])&(~a[3])&(a[2])&(a[1])&(a[0]);
assign y[24] = (a[4])&(a[3])&(~a[2])&(~a[1])&(~a[0]);
assign y[25] = (a[4])&(a[3])&(~a[2])&(~a[1])&(a[0]);
assign y[26] = (a[4])&(a[3])&(~a[2])&(a[1])&(~a[0]);
assign y[27] = (a[4])&(a[3])&(~a[2])&(a[1])&(a[0]);
assign y[28] = (a[4])&(a[3])&(a[2])&(~a[1])&(~a[0]);
assign y[29] = (a[4])&(a[3])&(a[2])&(~a[1])&(a[0]);
assign y[30] = (a[4])&(a[3])&(a[2])&(a[1])&(~a[0]);
assign y[31] = (a[4])&(a[3])&(a[2])&(a[1])&(a[0]);
endmodule
