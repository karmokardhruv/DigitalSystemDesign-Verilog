module and_gate(Y,a,b);
output Y; 
input a, b; 
and a_1(Y,a,b); 
endmodule
