module and_gate(a,b,Y);
input a,b;
output Y;
assign Y=a&b;
endmodule