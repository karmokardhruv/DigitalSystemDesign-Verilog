module xnor_gate(Y,a,b);
output Y;
input a, b;
xnor a_1(Y,a,b);
endmodule
